// This is a placeholder to disable IDE missing file warning.
// You should run sbt command first to generate this!

module $classname$ ();

endmodule
